module lcd_init (
    input wire clk,
    input wire rst_n,
    input wire spi_done,
    output reg spi_start,
    output reg [7:0] data_out
);

// Lógica para la inicialización de la pantalla LCD

endmodule
