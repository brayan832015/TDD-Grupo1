module spi_master (
    input wire clk,
    input wire rst_n,
    input wire start,
    input wire [7:0] data_in,
    output reg sck,
    output reg mosi,
    output reg cs_n,
    output reg done
);

// Lógica para el controlador SPI maestro

endmodule
