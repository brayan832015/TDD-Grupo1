module uart_rx (
    input wire clk,
    input wire rst_n,
    input wire rx,
    output reg [7:0] data_out,
    output reg ready
);

// Lógica de UART RX para recibir configuraciones de color desde la laptop

endmodule
