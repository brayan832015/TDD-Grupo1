module color_control (
    input wire clk,
    input wire rst_n,
    input wire [7:0] uart_data,
    input wire uart_ready,
    output reg [15:0] color_p1,
    output reg [15:0] color_p2
);

// Lógica para controlar las configuraciones de color

endmodule
